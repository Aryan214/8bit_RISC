module RISC_2Stage (
    input wire clk,
    input wire rst
);
    Datapath dp (.clk(clk), .rst(rst));
endmodule
